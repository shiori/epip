/// =============================================================================
///                         FILE DETAILS
/// Project          : IP4
/// Author           : Andy Chen
/// File             : ip4_rtl_bb.sv
/// Title            : ip4 building block
/// Version          : 0.1
/// Last modified    : Feb 21 2011
/// =============================================================================
///Log:
///Created by Andy Chen on Feb 21 2011

`ifdef IP4_ASIC_MODE


`else
`ifdef IP4_FPGA_MODE


`endif
`endif