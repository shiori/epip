
`include "ip4_tlm_if.svh"
`include "tlm_rec_pkg.sv"
`include "ip4_tlm_pkg.sv"

`undef IP4_TLM_PKG
`include "../misc/test_sys.sv"
`include "../misc/test.sv"
`include "../misc/top.sv"