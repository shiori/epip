
`include "ip4_tlm_if.svh"

`include "ip4_rtl_pkg.sv"
`include "ip4_tlm_pkg.sv"
`include "ip4_rtl_if.svh"

`include "ip4_rtl_bb.sv"
///`include "ip4_rtl_rfm.sv"
`include "ip4_rtl_spa.sv"
///`include "ip4_rtl_spu.sv"
///`include "ip4_rtl_ise.sv"
///`include "ip4_rtl_tlb.sv"
`include "ip4_rtl_dse.sv"
///`include "ip4_rtl_eif.sv"
///`include "ip4_rtl_ife.sv"
///`include "ip4_rtl_agent.sv"
`include "ip4_rtl_core.sv"

`include "../misc/top.sv"