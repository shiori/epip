/// =============================================================================
///                         FILE DETAILS
/// Project          : IP4
/// Author           : Andy Chen
/// File             : ip4_rtl_spa.sv
/// Title            : ip4 stream processor array
/// Version          : 0.1
/// Last modified    : Feb 7 2011
/// =============================================================================
///Log:
///Created by Andy Chen on Feb 7 2011

module ip4_rtl_spa(ip4_rtl_if.spa intf);


endmodule : ip4_rtl_spa

