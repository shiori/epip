
`ifndef IP4_RTL_SVH
`define IP4_RTL_SVH

`include "ip4_tlm_ts.svh"
import ip4_rtl_pkg::*;

`define IP4_ASIC_MODE
`define IP4_FPGA_MODE

`endif