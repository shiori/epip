
`include "ip4_tlm_if.svh"
`include "tlm_rec_pkg.sv"
`include "ip4_tlm_pkg.sv"
`include "../misc/top.sv"