
timeunit 1ns;
timeprecision 100ps;