
`ifdef IP4_RTL_PKG

`else

`ifndef IP4_RTL_SVH
`define IP4_RTL_SVH

`include "ip4_tlm_ts.svh"
import ip4_rtl_pkg::*;

`endif

`endif