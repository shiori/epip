
`include "ip4_tlm_if.svh"

`include "ip4_rtl_pkg.sv"
`include "ip4_tlm_pkg.sv"
`include "../misc/top.sv"